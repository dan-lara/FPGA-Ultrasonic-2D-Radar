library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TB_UART_Avalon_DUT is
end entity;

architecture Behavioral of TB_UART_Avalon_DUT is

    -- Signal
    signal clk        : std_logic := '0';
    signal Rst_n      : std_logic := '1';
    --signal load       : std_logic := '0';

    signal Read_n            : std_logic;
    signal ReadData          : std_logic_vector(31 downto 0);
    signal Write_n           : std_logic;
    signal WriteData         : std_logic_vector(31 downto 0) := (others => '0');

    signal Address           : std_logic_vector(1 downto 0) := (others => '0');


    --signal Tx_Data      : std_logic_vector(7 downto 0) := (others => '0');
    signal Uart_Tx      : std_logic;

    --signal Rx_Data      : std_logic_vector(7 downto 0);
    signal Uart_Rx            : std_logic := '1';
    
    -- Constants for clock generation
    constant CLK_PERIOD : time := 10 ns; -- 100 MHz clock

    -- Content
begin

    -- Instance of the entity under test
    DUT: entity work.IP_UART_Avalon
        port map (
            clk      => clk,
            Rst_n  => Rst_n,
            --Load     => load,

            Read_n    => Read_n,
            ReadData  => ReadData,
            Write_n   => Write_n,
            WriteData => WriteData,

            --Address   => Address,

            Uart_Tx  => Uart_Tx,
            --Tx_Data  => Tx_Data,
        
            Uart_Rx  => Uart_Rx
            --Rx_Data  => Rx_Data
        );
        
    -- Clock generation
    process
    begin
        while true loop
            clk <= '0';
            wait for CLK_PERIOD / 2;
            clk <= '1';
            wait for CLK_PERIOD / 2;
        end loop;
    end process;

    -- Test process
    process
    begin
        -- Initial reset
        Rst_n <= '0';
        wait for 50 ns;
        Rst_n <= '1';
        wait for 50 ns;
    
    -- Test Transmit
        -- D
        Read_n <= '1';
        Write_n <= '0';
        Address <= "01"; -- bits 31 et 30 
        WriteData <= "01000000000000000000000001000100";
        wait for CLK_PERIOD;
        Address <= "00";
        WriteData <= "00000000000000000000000000000001";--load <= '1';
        wait for 500*CLK_PERIOD;
        WriteData <= "00000000000000000000000000000000";--load <= '0';        
        wait for CLK_PERIOD;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";
        wait for 150 us;

        -- a
        Read_n <= '1';
        Write_n <= '0';
        Address <= "01";
        WriteData <= "01000000000000000000000001100001";
        wait for CLK_PERIOD;
        Address <= "00";
        WriteData <= "00000000000000000000000000000001";--load <= '1';
        wait for 500*CLK_PERIOD;
        WriteData <= "00000000000000000000000000000000";--load <= '0';        
        wait for CLK_PERIOD;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";
        WriteData <= "10000000000000000000000000000000";--load <= '0';
        wait for 150 us;

        --n
        Read_n <= '1';
        Write_n <= '0';
        Address <= "01";
        WriteData <= "01000000000000000000000001101110";
        wait for CLK_PERIOD;
        Address <= "00";
        WriteData <= "00000000000000000000000000000001";--load <= '1';
        wait for 500*CLK_PERIOD;
        WriteData <= "00000000000000000000000000000000";--load <= '0';        
        wait for CLK_PERIOD;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";
        WriteData <= "10000000000000000000000000000000";--load <= '0';
        wait for 150 us;

        --" "
        Read_n <= '1';
        Write_n <= '0';
        Address <= "01";
        WriteData <= "01000000000000000000000000100000";
        wait for CLK_PERIOD;
        Address <= "00";
        WriteData <= "00000000000000000000000000000001";--load <= '1';
        wait for 500*CLK_PERIOD;
        WriteData <= "00000000000000000000000000000000";--load <= '0';        
        wait for CLK_PERIOD;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";
        WriteData <= "10000000000000000000000000000000";--load <= '0';
        wait for 150 us;

        --L
        Read_n <= '1';
        Write_n <= '0';
        Address <= "01";
        WriteData <= "01000000000000000000000001001100";
        wait for CLK_PERIOD;
        Address <= "00";
        WriteData <= "00000000000000000000000000000001";--load <= '1';
        wait for 500*CLK_PERIOD;
        WriteData <= "00000000000000000000000000000000";--load <= '0';        
        wait for CLK_PERIOD;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";
        WriteData <= "10000000000000000000000000000000";--load <= '0';
        wait for 150 us;

        --"\n"
        Read_n <= '1';
        Write_n <= '0';
        Address <= "01";
        WriteData <= "01000000000000000000000000001010";
        wait for CLK_PERIOD;
        Address <= "00";
        WriteData <= "00000000000000000000000000000001";--load <= '1';
        wait for 500*CLK_PERIOD;
        WriteData <= "00000000000000000000000000000000";--load <= '0';        
        wait for CLK_PERIOD;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";
        WriteData <= "10000000000000000000000000000000";--load <= '0';
        wait for 150 us;

        -- Reseting
        Rst_n <= '0';
        wait for 70 us;

        Read_n <= '1';
        Write_n <= '0';
        Address <= "00";
        WriteData <= "00000000000000000000000000000001"; --load <= '1';
        wait for 30 us;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";

        wait for 50 us;

        Rst_n <= '1';
        Read_n <= '1';
        Write_n <= '0';
        Address <= "00";
        wait for 30 us;
        WriteData <= "00000000000000000000000000000000"; --load <= '0';
        wait for 30 us;
        Read_n <= '0';
        Write_n <= '1';
        Address <= "10";        
        WriteData <= "10000000000000000000000000000000";--load <= '0';

    -- Test Read
        wait for 160 us;
        Address <= "10";        
        WriteData <= "10000000000000000000000000000000";--load <= '0';

        -- Test case 0 : Read random data (ASCII '?')
        Uart_Rx <= '0';
        wait for 434*4*CLK_PERIOD;
        Uart_Rx <= '1';
        wait for 70 us;

        -- STOP_1 01001100 START_0
        Uart_Rx <= '0';
        wait for 434*CLK_PERIOD;
        wait for 434*CLK_PERIOD;
        wait for 434*CLK_PERIOD;
        Uart_Rx <= '1';
        wait for 434*CLK_PERIOD;
        wait for 434*CLK_PERIOD;
        Uart_Rx <= '0';
        wait for 434*CLK_PERIOD;
        wait for 434*CLK_PERIOD;
        Uart_Rx <= '1';
        wait for 434*CLK_PERIOD;
        Uart_Rx <= '0';
        wait for 434*CLK_PERIOD;
        Uart_Rx <= '1';
        wait for 30 us;


        -- End simulation
        wait;
    end process;

end architecture;