// Computer_System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Computer_System (
		inout  wire [15:0] arduino_gpio_export,        //         arduino_gpio.export
		output wire        arduino_reset_n_export,     //      arduino_reset_n.export
		output wire [31:0] hex3_hex0_export,           //            hex3_hex0.export
		output wire [15:0] hex5_hex4_export,           //            hex5_hex4.export
		output wire [9:0]  leds_export,                //                 leds.export
		output wire        neopixel_out_commande,      //         neopixel_out.commande
		input  wire [1:0]  pushbuttons_export,         //          pushbuttons.export
		output wire [12:0] sdram_addr,                 //                sdram.addr
		output wire [1:0]  sdram_ba,                   //                     .ba
		output wire        sdram_cas_n,                //                     .cas_n
		output wire        sdram_cke,                  //                     .cke
		output wire        sdram_cs_n,                 //                     .cs_n
		inout  wire [15:0] sdram_dq,                   //                     .dq
		output wire [1:0]  sdram_dqm,                  //                     .dqm
		output wire        sdram_ras_n,                //                     .ras_n
		output wire        sdram_we_n,                 //                     .we_n
		output wire        sdram_clk_clk,              //            sdram_clk.clk
		output wire        servo_out_commande,         //            servo_out.commande
		input  wire [9:0]  slider_switches_export,     //      slider_switches.export
		input  wire        system_pll_ref_clk_clk,     //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset, // system_pll_ref_reset.reset
		output wire [9:0]  telemetre_out_dist_cm,      //        telemetre_out.dist_cm
		input  wire        telemetre_out_echo,         //                     .echo
		output wire        telemetre_out_trig,         //                     .trig
		input  wire        uart_out_commande_rx,       //             uart_out.commande_rx
		output wire        uart_out_commande_tx,       //                     .commande_tx
		output wire        vga_CLK,                    //                  vga.CLK
		output wire        vga_HS,                     //                     .HS
		output wire        vga_VS,                     //                     .VS
		output wire        vga_BLANK,                  //                     .BLANK
		output wire        vga_SYNC,                   //                     .SYNC
		output wire [3:0]  vga_R,                      //                     .R
		output wire [3:0]  vga_G,                      //                     .G
		output wire [3:0]  vga_B,                      //                     .B
		input  wire        video_pll_ref_clk_clk,      //    video_pll_ref_clk.clk
		input  wire        video_pll_ref_reset_reset   //  video_pll_ref_reset.reset
	);

	wire         system_pll_sys_clk_clk;                                                   // System_PLL:sys_clk_clk -> [Arduino_GPIO:clk, Arduino_Reset_N:clk, HEX3_HEX0:clk, HEX5_HEX4:clk, Interval_Timer:clk, Interval_Timer_2:clk, JTAG_UART:clk, JTAG_to_FPGA_Bridge:clk_clk, LEDs:clk, Nios2:clk, Onchip_SRAM:clk, Pushbuttons:clk, SDRAM:clk, Slider_Switches:clk, SysID:clock, VGA_Subsystem:sys_clk_clk, irq_mapper:clk, mm_interconnect_0:System_PLL_sys_clk_clk, neopixel_0:clk, rst_controller:clk, rst_controller_001:clk, servo_0:clk, telemetre_0:clk, uart_0:clk]
	wire         video_pll_vga_clk_clk;                                                    // Video_PLL:vga_clk_clk -> VGA_Subsystem:vga_clk_clk
	wire         system_pll_reset_source_reset;                                            // System_PLL:reset_source_reset -> [JTAG_to_FPGA_Bridge:clk_reset_reset, VGA_Subsystem:sys_reset_reset_n, rst_controller:reset_in0, rst_controller_001:reset_in1]
	wire         video_pll_reset_source_reset;                                             // Video_PLL:reset_source_reset -> VGA_Subsystem:vga_reset_reset_n
	wire         nios2_custom_instruction_master_readra;                                   // Nios2:D_ci_readra -> Nios2_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_a;                                        // Nios2:D_ci_a -> Nios2_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_b;                                        // Nios2:D_ci_b -> Nios2_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_custom_instruction_master_c;                                        // Nios2:D_ci_c -> Nios2_custom_instruction_master_translator:ci_slave_c
	wire         nios2_custom_instruction_master_readrb;                                   // Nios2:D_ci_readrb -> Nios2_custom_instruction_master_translator:ci_slave_readrb
	wire         nios2_custom_instruction_master_clk;                                      // Nios2:E_ci_multi_clock -> Nios2_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_custom_instruction_master_ipending;                                 // Nios2:W_ci_ipending -> Nios2_custom_instruction_master_translator:ci_slave_ipending
	wire         nios2_custom_instruction_master_start;                                    // Nios2:E_ci_multi_start -> Nios2_custom_instruction_master_translator:ci_slave_multi_start
	wire         nios2_custom_instruction_master_reset_req;                                // Nios2:E_ci_multi_reset_req -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_custom_instruction_master_done;                                     // Nios2_custom_instruction_master_translator:ci_slave_multi_done -> Nios2:E_ci_multi_done
	wire   [7:0] nios2_custom_instruction_master_n;                                        // Nios2:D_ci_n -> Nios2_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_result;                                   // Nios2_custom_instruction_master_translator:ci_slave_result -> Nios2:E_ci_result
	wire         nios2_custom_instruction_master_estatus;                                  // Nios2:W_ci_estatus -> Nios2_custom_instruction_master_translator:ci_slave_estatus
	wire         nios2_custom_instruction_master_clk_en;                                   // Nios2:E_ci_multi_clk_en -> Nios2_custom_instruction_master_translator:ci_slave_multi_clken
	wire  [31:0] nios2_custom_instruction_master_datab;                                    // Nios2:E_ci_datab -> Nios2_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_dataa;                                    // Nios2:E_ci_dataa -> Nios2_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_custom_instruction_master_reset;                                    // Nios2:E_ci_multi_reset -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_custom_instruction_master_writerc;                                  // Nios2:D_ci_writerc -> Nios2_custom_instruction_master_translator:ci_slave_writerc
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readra;        // Nios2_custom_instruction_master_translator:multi_ci_master_readra -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_a;             // Nios2_custom_instruction_master_translator:multi_ci_master_a -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_b;             // Nios2_custom_instruction_master_translator:multi_ci_master_b -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk;           // Nios2_custom_instruction_master_translator:multi_ci_master_clk -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readrb;        // Nios2_custom_instruction_master_translator:multi_ci_master_readrb -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_c;             // Nios2_custom_instruction_master_translator:multi_ci_master_c -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_custom_instruction_master_translator_multi_ci_master_start;         // Nios2_custom_instruction_master_translator:multi_ci_master_start -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset_req;     // Nios2_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_custom_instruction_master_translator_multi_ci_master_done;          // Nios2_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios2_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_custom_instruction_master_translator_multi_ci_master_n;             // Nios2_custom_instruction_master_translator:multi_ci_master_n -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_result;        // Nios2_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios2_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk_en;        // Nios2_custom_instruction_master_translator:multi_ci_master_clken -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_datab;         // Nios2_custom_instruction_master_translator:multi_ci_master_datab -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_dataa;         // Nios2_custom_instruction_master_translator:multi_ci_master_dataa -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset;         // Nios2_custom_instruction_master_translator:multi_ci_master_reset -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_custom_instruction_master_translator_multi_ci_master_writerc;       // Nios2_custom_instruction_master_translator:multi_ci_master_writerc -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readra;         // Nios2_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_a;              // Nios2_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_b;              // Nios2_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb;         // Nios2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_c;              // Nios2_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk;            // Nios2_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending;       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_start;          // Nios2_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req;      // Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_done;           // Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_n;              // Nios2_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_result;         // Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus;        // Nios2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en;         // Nios2_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_datab;          // Nios2_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa;          // Nios2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset;          // Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc;        // Nios2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_result; // Nios2_Floating_Point:result -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk;    // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_Floating_Point:clk
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en; // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_Floating_Point:clk_en
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab;  // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_Floating_Point:datab
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa;  // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_Floating_Point:dataa
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_start;  // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_Floating_Point:start
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset;  // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_Floating_Point:reset
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_done;   // Nios2_Floating_Point:done -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [1:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_n;      // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_Floating_Point:n
	wire  [31:0] nios2_data_master_readdata;                                               // mm_interconnect_0:Nios2_data_master_readdata -> Nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                            // mm_interconnect_0:Nios2_data_master_waitrequest -> Nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                            // Nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_data_master_debugaccess
	wire  [31:0] nios2_data_master_address;                                                // Nios2:d_address -> mm_interconnect_0:Nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                             // Nios2:d_byteenable -> mm_interconnect_0:Nios2_data_master_byteenable
	wire         nios2_data_master_read;                                                   // Nios2:d_read -> mm_interconnect_0:Nios2_data_master_read
	wire         nios2_data_master_write;                                                  // Nios2:d_write -> mm_interconnect_0:Nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                              // Nios2:d_writedata -> mm_interconnect_0:Nios2_data_master_writedata
	wire  [31:0] jtag_to_fpga_bridge_master_readdata;                                      // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	wire         jtag_to_fpga_bridge_master_waitrequest;                                   // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	wire  [31:0] jtag_to_fpga_bridge_master_address;                                       // JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_address
	wire         jtag_to_fpga_bridge_master_read;                                          // JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_read
	wire   [3:0] jtag_to_fpga_bridge_master_byteenable;                                    // JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_byteenable
	wire         jtag_to_fpga_bridge_master_readdatavalid;                                 // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	wire         jtag_to_fpga_bridge_master_write;                                         // JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_write
	wire  [31:0] jtag_to_fpga_bridge_master_writedata;                                     // JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                                        // mm_interconnect_0:Nios2_instruction_master_readdata -> Nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                                     // mm_interconnect_0:Nios2_instruction_master_waitrequest -> Nios2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                                         // Nios2:i_address -> mm_interconnect_0:Nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                            // Nios2:i_read -> mm_interconnect_0:Nios2_instruction_master_read
	wire         vga_subsystem_pixel_dma_master_waitrequest;                               // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_waitrequest -> VGA_Subsystem:pixel_dma_master_waitrequest
	wire  [15:0] vga_subsystem_pixel_dma_master_readdata;                                  // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdata -> VGA_Subsystem:pixel_dma_master_readdata
	wire  [31:0] vga_subsystem_pixel_dma_master_address;                                   // VGA_Subsystem:pixel_dma_master_address -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_address
	wire         vga_subsystem_pixel_dma_master_read;                                      // VGA_Subsystem:pixel_dma_master_read -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_read
	wire         vga_subsystem_pixel_dma_master_readdatavalid;                             // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdatavalid -> VGA_Subsystem:pixel_dma_master_readdatavalid
	wire         vga_subsystem_pixel_dma_master_lock;                                      // VGA_Subsystem:pixel_dma_master_lock -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_lock
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                 // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                   // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                    // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                      // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                  // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire         mm_interconnect_0_telemetre_0_avalon_slave_0_chipselect;                  // mm_interconnect_0:telemetre_0_avalon_slave_0_chipselect -> telemetre_0:chipselect
	wire  [31:0] mm_interconnect_0_telemetre_0_avalon_slave_0_readdata;                    // telemetre_0:readdata -> mm_interconnect_0:telemetre_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_telemetre_0_avalon_slave_0_read;                        // mm_interconnect_0:telemetre_0_avalon_slave_0_read -> telemetre_0:Read_n
	wire         mm_interconnect_0_servo_0_avalon_slave_0_chipselect;                      // mm_interconnect_0:servo_0_avalon_slave_0_chipselect -> servo_0:chipselect
	wire         mm_interconnect_0_servo_0_avalon_slave_0_write;                           // mm_interconnect_0:servo_0_avalon_slave_0_write -> servo_0:write_n
	wire  [31:0] mm_interconnect_0_servo_0_avalon_slave_0_writedata;                       // mm_interconnect_0:servo_0_avalon_slave_0_writedata -> servo_0:WriteData
	wire         mm_interconnect_0_neopixel_0_avalon_slave_0_chipselect;                   // mm_interconnect_0:neopixel_0_avalon_slave_0_chipselect -> neopixel_0:chipselect
	wire         mm_interconnect_0_neopixel_0_avalon_slave_0_write;                        // mm_interconnect_0:neopixel_0_avalon_slave_0_write -> neopixel_0:write_n
	wire  [31:0] mm_interconnect_0_neopixel_0_avalon_slave_0_writedata;                    // mm_interconnect_0:neopixel_0_avalon_slave_0_writedata -> neopixel_0:WriteData
	wire  [31:0] mm_interconnect_0_uart_0_avalon_slave_0_readdata;                         // uart_0:ReadData -> mm_interconnect_0:uart_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_uart_0_avalon_slave_0_read;                             // mm_interconnect_0:uart_0_avalon_slave_0_read -> uart_0:Read_n
	wire         mm_interconnect_0_uart_0_avalon_slave_0_write;                            // mm_interconnect_0:uart_0_avalon_slave_0_write -> uart_0:Write_n
	wire  [31:0] mm_interconnect_0_uart_0_avalon_slave_0_writedata;                        // mm_interconnect_0:uart_0_avalon_slave_0_writedata -> uart_0:WriteData
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata;       // VGA_Subsystem:char_buffer_control_slave_readdata -> mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address;        // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_address -> VGA_Subsystem:char_buffer_control_slave_address
	wire         mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read;           // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_read -> VGA_Subsystem:char_buffer_control_slave_read
	wire   [3:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable;     // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_byteenable -> VGA_Subsystem:char_buffer_control_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write;          // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_write -> VGA_Subsystem:char_buffer_control_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata;      // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_writedata -> VGA_Subsystem:char_buffer_control_slave_writedata
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect;             // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_chipselect -> VGA_Subsystem:char_buffer_slave_chipselect
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata;               // VGA_Subsystem:char_buffer_slave_readdata -> mm_interconnect_0:VGA_Subsystem_char_buffer_slave_readdata
	wire  [10:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_address;                // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_address -> VGA_Subsystem:char_buffer_slave_address
	wire   [3:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable;             // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_byteenable -> VGA_Subsystem:char_buffer_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_write;                  // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_write -> VGA_Subsystem:char_buffer_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata;              // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_writedata -> VGA_Subsystem:char_buffer_slave_writedata
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_clken;                  // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_clken -> VGA_Subsystem:char_buffer_slave_clken
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                           // SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                            // mm_interconnect_0:SysID_control_slave_address -> SysID:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                         // Nios2:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;                      // Nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;                      // mm_interconnect_0:Nios2_debug_mem_slave_debugaccess -> Nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                          // mm_interconnect_0:Nios2_debug_mem_slave_address -> Nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                             // mm_interconnect_0:Nios2_debug_mem_slave_read -> Nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                       // mm_interconnect_0:Nios2_debug_mem_slave_byteenable -> Nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                            // mm_interconnect_0:Nios2_debug_mem_slave_write -> Nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                        // mm_interconnect_0:Nios2_debug_mem_slave_writedata -> Nios2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata;         // VGA_Subsystem:pixel_dma_control_slave_readdata -> mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address;          // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_address -> VGA_Subsystem:pixel_dma_control_slave_address
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read;             // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_read -> VGA_Subsystem:pixel_dma_control_slave_read
	wire   [3:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable;       // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_byteenable -> VGA_Subsystem:pixel_dma_control_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write;            // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_write -> VGA_Subsystem:pixel_dma_control_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata;        // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_writedata -> VGA_Subsystem:pixel_dma_control_slave_writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_rgb_slave_readdata;                       // VGA_Subsystem:rgb_slave_readdata -> mm_interconnect_0:VGA_Subsystem_rgb_slave_readdata
	wire         mm_interconnect_0_vga_subsystem_rgb_slave_read;                           // mm_interconnect_0:VGA_Subsystem_rgb_slave_read -> VGA_Subsystem:rgb_slave_read
	wire         mm_interconnect_0_sdram_s1_chipselect;                                    // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                      // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                   // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                       // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                          // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                    // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                 // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                         // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                     // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_onchip_sram_s1_chipselect;                              // mm_interconnect_0:Onchip_SRAM_s1_chipselect -> Onchip_SRAM:chipselect
	wire  [31:0] mm_interconnect_0_onchip_sram_s1_readdata;                                // Onchip_SRAM:readdata -> mm_interconnect_0:Onchip_SRAM_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_sram_s1_address;                                 // mm_interconnect_0:Onchip_SRAM_s1_address -> Onchip_SRAM:address
	wire   [3:0] mm_interconnect_0_onchip_sram_s1_byteenable;                              // mm_interconnect_0:Onchip_SRAM_s1_byteenable -> Onchip_SRAM:byteenable
	wire         mm_interconnect_0_onchip_sram_s1_write;                                   // mm_interconnect_0:Onchip_SRAM_s1_write -> Onchip_SRAM:write
	wire  [31:0] mm_interconnect_0_onchip_sram_s1_writedata;                               // mm_interconnect_0:Onchip_SRAM_s1_writedata -> Onchip_SRAM:writedata
	wire         mm_interconnect_0_onchip_sram_s1_clken;                                   // mm_interconnect_0:Onchip_SRAM_s1_clken -> Onchip_SRAM:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                                     // mm_interconnect_0:LEDs_s1_chipselect -> LEDs:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                       // LEDs:readdata -> mm_interconnect_0:LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                        // mm_interconnect_0:LEDs_s1_address -> LEDs:address
	wire         mm_interconnect_0_leds_s1_write;                                          // mm_interconnect_0:LEDs_s1_write -> LEDs:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                      // mm_interconnect_0:LEDs_s1_writedata -> LEDs:writedata
	wire         mm_interconnect_0_hex3_hex0_s1_chipselect;                                // mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_readdata;                                  // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_hex0_s1_address;                                   // mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_s1_write;                                     // mm_interconnect_0:HEX3_HEX0_s1_write -> HEX3_HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_writedata;                                 // mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	wire         mm_interconnect_0_hex5_hex4_s1_chipselect;                                // mm_interconnect_0:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_readdata;                                  // HEX5_HEX4:readdata -> mm_interconnect_0:HEX5_HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_hex4_s1_address;                                   // mm_interconnect_0:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	wire         mm_interconnect_0_hex5_hex4_s1_write;                                     // mm_interconnect_0:HEX5_HEX4_s1_write -> HEX5_HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_writedata;                                 // mm_interconnect_0:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	wire  [31:0] mm_interconnect_0_slider_switches_s1_readdata;                            // Slider_Switches:readdata -> mm_interconnect_0:Slider_Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_slider_switches_s1_address;                             // mm_interconnect_0:Slider_Switches_s1_address -> Slider_Switches:address
	wire         mm_interconnect_0_pushbuttons_s1_chipselect;                              // mm_interconnect_0:Pushbuttons_s1_chipselect -> Pushbuttons:chipselect
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_readdata;                                // Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_s1_address;                                 // mm_interconnect_0:Pushbuttons_s1_address -> Pushbuttons:address
	wire         mm_interconnect_0_pushbuttons_s1_write;                                   // mm_interconnect_0:Pushbuttons_s1_write -> Pushbuttons:write_n
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_writedata;                               // mm_interconnect_0:Pushbuttons_s1_writedata -> Pushbuttons:writedata
	wire         mm_interconnect_0_arduino_gpio_s1_chipselect;                             // mm_interconnect_0:Arduino_GPIO_s1_chipselect -> Arduino_GPIO:chipselect
	wire  [31:0] mm_interconnect_0_arduino_gpio_s1_readdata;                               // Arduino_GPIO:readdata -> mm_interconnect_0:Arduino_GPIO_s1_readdata
	wire   [1:0] mm_interconnect_0_arduino_gpio_s1_address;                                // mm_interconnect_0:Arduino_GPIO_s1_address -> Arduino_GPIO:address
	wire         mm_interconnect_0_arduino_gpio_s1_write;                                  // mm_interconnect_0:Arduino_GPIO_s1_write -> Arduino_GPIO:write_n
	wire  [31:0] mm_interconnect_0_arduino_gpio_s1_writedata;                              // mm_interconnect_0:Arduino_GPIO_s1_writedata -> Arduino_GPIO:writedata
	wire         mm_interconnect_0_arduino_reset_n_s1_chipselect;                          // mm_interconnect_0:Arduino_Reset_N_s1_chipselect -> Arduino_Reset_N:chipselect
	wire  [31:0] mm_interconnect_0_arduino_reset_n_s1_readdata;                            // Arduino_Reset_N:readdata -> mm_interconnect_0:Arduino_Reset_N_s1_readdata
	wire   [1:0] mm_interconnect_0_arduino_reset_n_s1_address;                             // mm_interconnect_0:Arduino_Reset_N_s1_address -> Arduino_Reset_N:address
	wire         mm_interconnect_0_arduino_reset_n_s1_write;                               // mm_interconnect_0:Arduino_Reset_N_s1_write -> Arduino_Reset_N:write_n
	wire  [31:0] mm_interconnect_0_arduino_reset_n_s1_writedata;                           // mm_interconnect_0:Arduino_Reset_N_s1_writedata -> Arduino_Reset_N:writedata
	wire         mm_interconnect_0_interval_timer_s1_chipselect;                           // mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_s1_readdata;                             // Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_s1_address;                              // mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	wire         mm_interconnect_0_interval_timer_s1_write;                                // mm_interconnect_0:Interval_Timer_s1_write -> Interval_Timer:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_s1_writedata;                            // mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	wire         mm_interconnect_0_interval_timer_2_s1_chipselect;                         // mm_interconnect_0:Interval_Timer_2_s1_chipselect -> Interval_Timer_2:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_2_s1_readdata;                           // Interval_Timer_2:readdata -> mm_interconnect_0:Interval_Timer_2_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_2_s1_address;                            // mm_interconnect_0:Interval_Timer_2_s1_address -> Interval_Timer_2:address
	wire         mm_interconnect_0_interval_timer_2_s1_write;                              // mm_interconnect_0:Interval_Timer_2_s1_write -> Interval_Timer_2:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_2_s1_writedata;                          // mm_interconnect_0:Interval_Timer_2_s1_writedata -> Interval_Timer_2:writedata
	wire         mm_interconnect_0_onchip_sram_s2_chipselect;                              // mm_interconnect_0:Onchip_SRAM_s2_chipselect -> Onchip_SRAM:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_sram_s2_readdata;                                // Onchip_SRAM:readdata2 -> mm_interconnect_0:Onchip_SRAM_s2_readdata
	wire  [13:0] mm_interconnect_0_onchip_sram_s2_address;                                 // mm_interconnect_0:Onchip_SRAM_s2_address -> Onchip_SRAM:address2
	wire   [3:0] mm_interconnect_0_onchip_sram_s2_byteenable;                              // mm_interconnect_0:Onchip_SRAM_s2_byteenable -> Onchip_SRAM:byteenable2
	wire         mm_interconnect_0_onchip_sram_s2_write;                                   // mm_interconnect_0:Onchip_SRAM_s2_write -> Onchip_SRAM:write2
	wire  [31:0] mm_interconnect_0_onchip_sram_s2_writedata;                               // mm_interconnect_0:Onchip_SRAM_s2_writedata -> Onchip_SRAM:writedata2
	wire         mm_interconnect_0_onchip_sram_s2_clken;                                   // mm_interconnect_0:Onchip_SRAM_s2_clken -> Onchip_SRAM:clken2
	wire         irq_mapper_receiver0_irq;                                                 // Pushbuttons:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                 // Arduino_GPIO:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                 // JTAG_UART:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                 // Interval_Timer:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                 // Interval_Timer_2:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_irq_irq;                                                            // irq_mapper:sender_irq -> Nios2:irq
	wire         rst_controller_reset_out_reset;                                           // rst_controller:reset_out -> [Arduino_GPIO:reset_n, Arduino_Reset_N:reset_n, HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, Interval_Timer:reset_n, Interval_Timer_2:reset_n, JTAG_UART:rst_n, LEDs:reset_n, Onchip_SRAM:reset, Pushbuttons:reset_n, SDRAM:reset_n, Slider_Switches:reset_n, SysID:reset_n, mm_interconnect_0:JTAG_UART_reset_reset_bridge_in_reset_reset, mm_interconnect_0:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, neopixel_0:Rst_n, rst_translator:in_reset, servo_0:reset_n, telemetre_0:Rst_n, uart_0:Rst_n]
	wire         rst_controller_reset_out_reset_req;                                       // rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                       // rst_controller_001:reset_out -> [Nios2:reset_n, irq_mapper:reset, mm_interconnect_0:Nios2_reset_reset_bridge_in_reset_reset]
	wire         nios2_debug_reset_request_reset;                                          // Nios2:debug_reset_request -> rst_controller_001:reset_in0

	Computer_System_Arduino_GPIO arduino_gpio (
		.clk        (system_pll_sys_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_arduino_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_arduino_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_arduino_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_arduino_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_arduino_gpio_s1_readdata),   //                    .readdata
		.bidir_port (arduino_gpio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                      //                 irq.irq
	);

	Computer_System_Arduino_Reset_N arduino_reset_n (
		.clk        (system_pll_sys_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_arduino_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_arduino_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_arduino_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_arduino_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_arduino_reset_n_s1_readdata),   //                    .readdata
		.out_port   (arduino_reset_n_export)                           // external_connection.export
	);

	Computer_System_HEX3_HEX0 hex3_hex0 (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex3_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex3_hex0_export)                           // external_connection.export
	);

	Computer_System_HEX5_HEX4 hex5_hex4 (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex5_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex5_hex4_export)                           // external_connection.export
	);

	Computer_System_Interval_Timer interval_timer (
		.clk        (system_pll_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                        //   irq.irq
	);

	Computer_System_Interval_Timer interval_timer_2 (
		.clk        (system_pll_sys_clk_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_2_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                          //   irq.irq
	);

	Computer_System_JTAG_UART jtag_uart (
		.clk            (system_pll_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	Computer_System_JTAG_to_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_fpga_bridge (
		.clk_clk              (system_pll_sys_clk_clk),                   //          clk.clk
		.clk_reset_reset      (system_pll_reset_source_reset),            //    clk_reset.reset
		.master_address       (jtag_to_fpga_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_fpga_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_fpga_bridge_master_read),          //             .read
		.master_write         (jtag_to_fpga_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_fpga_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_fpga_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_fpga_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_fpga_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	Computer_System_LEDs leds (
		.clk        (system_pll_sys_clk_clk),               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	Computer_System_Nios2 nios2 (
		.clk                                 (system_pll_sys_clk_clk),                              //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_multi_done                     (nios2_custom_instruction_master_done),                // custom_instruction_master.done
		.E_ci_multi_clk_en                   (nios2_custom_instruction_master_clk_en),              //                          .clk_en
		.E_ci_multi_start                    (nios2_custom_instruction_master_start),               //                          .start
		.E_ci_result                         (nios2_custom_instruction_master_result),              //                          .result
		.D_ci_a                              (nios2_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (nios2_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (nios2_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (nios2_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (nios2_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (nios2_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (nios2_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (nios2_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (nios2_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (nios2_custom_instruction_master_clk),                 //                          .clk
		.E_ci_multi_reset                    (nios2_custom_instruction_master_reset),               //                          .reset
		.E_ci_multi_reset_req                (nios2_custom_instruction_master_reset_req),           //                          .reset_req
		.W_ci_estatus                        (nios2_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (nios2_custom_instruction_master_ipending)             //                          .ipending
	);

	fpoint_wrapper #(
		.useDivider (1)
	) nios2_floating_point (
		.clk    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // s1.clk
		.clk_en (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //   .clk_en
		.dataa  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //   .dataa
		.datab  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //   .datab
		.n      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //   .n
		.reset  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //   .reset
		.start  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //   .start
		.done   (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //   .done
		.result (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result)  //   .result
	);

	Computer_System_Onchip_SRAM onchip_sram (
		.address     (mm_interconnect_0_onchip_sram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_sram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_sram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_sram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_sram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_sram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_sram_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_sram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_sram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_sram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_sram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_sram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_sram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_sram_s2_byteenable), //       .byteenable
		.clk         (system_pll_sys_clk_clk),                      //   clk1.clk
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	Computer_System_Pushbuttons pushbuttons (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pushbuttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbuttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbuttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbuttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbuttons_s1_readdata),   //                    .readdata
		.in_port    (pushbuttons_export),                          // external_connection.export
		.irq        (irq_mapper_receiver0_irq)                     //                 irq.irq
	);

	Computer_System_SDRAM sdram (
		.clk            (system_pll_sys_clk_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	Computer_System_Slider_Switches slider_switches (
		.clk      (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_slider_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_slider_switches_s1_readdata), //                    .readdata
		.in_port  (slider_switches_export)                         // external_connection.export
	);

	Computer_System_SysID sysid (
		.clock    (system_pll_sys_clk_clk),                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_VGA_Subsystem vga_subsystem (
		.char_buffer_control_slave_address    (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address),    // char_buffer_control_slave.address
		.char_buffer_control_slave_byteenable (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable), //                          .byteenable
		.char_buffer_control_slave_read       (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read),       //                          .read
		.char_buffer_control_slave_write      (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write),      //                          .write
		.char_buffer_control_slave_writedata  (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata),  //                          .writedata
		.char_buffer_control_slave_readdata   (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata),   //                          .readdata
		.char_buffer_slave_address            (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),            //         char_buffer_slave.address
		.char_buffer_slave_clken              (mm_interconnect_0_vga_subsystem_char_buffer_slave_clken),              //                          .clken
		.char_buffer_slave_chipselect         (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect),         //                          .chipselect
		.char_buffer_slave_write              (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),              //                          .write
		.char_buffer_slave_readdata           (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),           //                          .readdata
		.char_buffer_slave_writedata          (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),          //                          .writedata
		.char_buffer_slave_byteenable         (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),         //                          .byteenable
		.pixel_dma_control_slave_address      (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),      //   pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable   (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable),   //                          .byteenable
		.pixel_dma_control_slave_read         (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),         //                          .read
		.pixel_dma_control_slave_write        (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),        //                          .write
		.pixel_dma_control_slave_writedata    (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),    //                          .writedata
		.pixel_dma_control_slave_readdata     (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),     //                          .readdata
		.pixel_dma_master_address             (vga_subsystem_pixel_dma_master_address),                               //          pixel_dma_master.address
		.pixel_dma_master_waitrequest         (vga_subsystem_pixel_dma_master_waitrequest),                           //                          .waitrequest
		.pixel_dma_master_lock                (vga_subsystem_pixel_dma_master_lock),                                  //                          .lock
		.pixel_dma_master_read                (vga_subsystem_pixel_dma_master_read),                                  //                          .read
		.pixel_dma_master_readdata            (vga_subsystem_pixel_dma_master_readdata),                              //                          .readdata
		.pixel_dma_master_readdatavalid       (vga_subsystem_pixel_dma_master_readdatavalid),                         //                          .readdatavalid
		.rgb_slave_read                       (mm_interconnect_0_vga_subsystem_rgb_slave_read),                       //                 rgb_slave.read
		.rgb_slave_readdata                   (mm_interconnect_0_vga_subsystem_rgb_slave_readdata),                   //                          .readdata
		.sys_clk_clk                          (system_pll_sys_clk_clk),                                               //                   sys_clk.clk
		.sys_reset_reset_n                    (~system_pll_reset_source_reset),                                       //                 sys_reset.reset_n
		.vga_CLK                              (vga_CLK),                                                              //                       vga.CLK
		.vga_HS                               (vga_HS),                                                               //                          .HS
		.vga_VS                               (vga_VS),                                                               //                          .VS
		.vga_BLANK                            (vga_BLANK),                                                            //                          .BLANK
		.vga_SYNC                             (vga_SYNC),                                                             //                          .SYNC
		.vga_R                                (vga_R),                                                                //                          .R
		.vga_G                                (vga_G),                                                                //                          .G
		.vga_B                                (vga_B),                                                                //                          .B
		.vga_clk_clk                          (video_pll_vga_clk_clk),                                                //                   vga_clk.clk
		.vga_reset_reset_n                    (~video_pll_reset_source_reset)                                         //                 vga_reset.reset_n
	);

	Computer_System_Video_PLL video_pll (
		.ref_clk_clk        (video_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (video_pll_ref_reset_reset),    //    ref_reset.reset
		.vga_clk_clk        (video_pll_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_reset_source_reset)  // reset_source.reset
	);

	IP_NeoPixel_Avalon neopixel_0 (
		.clk        (system_pll_sys_clk_clk),                                 //          clock.clk
		.chipselect (mm_interconnect_0_neopixel_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.write_n    (~mm_interconnect_0_neopixel_0_avalon_slave_0_write),     //               .write_n
		.WriteData  (mm_interconnect_0_neopixel_0_avalon_slave_0_writedata),  //               .writedata
		.Rst_n      (~rst_controller_reset_out_reset),                        //     reset_sink.reset_n
		.commande   (neopixel_out_commande)                                   //    conduit_end.commande
	);

	IP_Servo_Avalon servo_0 (
		.clk        (system_pll_sys_clk_clk),                              //          clock.clk
		.chipselect (mm_interconnect_0_servo_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.write_n    (~mm_interconnect_0_servo_0_avalon_slave_0_write),     //               .write_n
		.WriteData  (mm_interconnect_0_servo_0_avalon_slave_0_writedata),  //               .writedata
		.commande   (servo_out_commande),                                  //    conduit_end.commande
		.reset_n    (~rst_controller_reset_out_reset)                      //     reset_sink.reset_n
	);

	IP_Telemetre_Avalon telemetre_0 (
		.clk        (system_pll_sys_clk_clk),                                  //          clock.clk
		.chipselect (mm_interconnect_0_telemetre_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.Read_n     (~mm_interconnect_0_telemetre_0_avalon_slave_0_read),      //               .read_n
		.readdata   (mm_interconnect_0_telemetre_0_avalon_slave_0_readdata),   //               .readdata
		.Dist_cm    (telemetre_out_dist_cm),                                   //    conduit_end.dist_cm
		.echo       (telemetre_out_echo),                                      //               .echo
		.trig       (telemetre_out_trig),                                      //               .trig
		.Rst_n      (~rst_controller_reset_out_reset)                          //     reset_sink.reset_n
	);

	IP_UART_Avalon uart_0 (
		.clk       (system_pll_sys_clk_clk),                            //          clock.clk
		.Read_n    (~mm_interconnect_0_uart_0_avalon_slave_0_read),     // avalon_slave_0.read_n
		.ReadData  (mm_interconnect_0_uart_0_avalon_slave_0_readdata),  //               .readdata
		.Write_n   (~mm_interconnect_0_uart_0_avalon_slave_0_write),    //               .write_n
		.WriteData (mm_interconnect_0_uart_0_avalon_slave_0_writedata), //               .writedata
		.Uart_Rx   (uart_out_commande_rx),                              //    conduit_end.commande_rx
		.Uart_Tx   (uart_out_commande_tx),                              //               .commande_tx
		.Rst_n     (~rst_controller_reset_out_reset)                    //     reset_sink.reset_n
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (nios2_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (nios2_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (nios2_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (nios2_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (nios2_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (nios2_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (nios2_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (nios2_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (nios2_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (nios2_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (nios2_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (nios2_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (),                                                                     //  comb_ci_master.dataa
		.comb_ci_master_datab      (),                                                                     //                .datab
		.comb_ci_master_result     (),                                                                     //                .result
		.comb_ci_master_n          (),                                                                     //                .n
		.comb_ci_master_readra     (),                                                                     //                .readra
		.comb_ci_master_readrb     (),                                                                     //                .readrb
		.comb_ci_master_writerc    (),                                                                     //                .writerc
		.comb_ci_master_a          (),                                                                     //                .a
		.comb_ci_master_b          (),                                                                     //                .b
		.comb_ci_master_c          (),                                                                     //                .c
		.comb_ci_master_ipending   (),                                                                     //                .ipending
		.comb_ci_master_estatus    (),                                                                     //                .estatus
		.multi_ci_master_clk       (nios2_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_multi_result     (),                                                                     //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                          //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                 //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                 //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                 //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                             //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                             //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                              //     (terminated)
	);

	Computer_System_Nios2_custom_instruction_master_multi_xconnect nios2_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (nios2_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_reset_req ()                                                                          // (terminated)
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.System_PLL_sys_clk_clk                                    (system_pll_sys_clk_clk),                                               //                                  System_PLL_sys_clk.clk
		.JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                       // JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
		.JTAG_UART_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                       //               JTAG_UART_reset_reset_bridge_in_reset.reset
		.Nios2_reset_reset_bridge_in_reset_reset                   (rst_controller_001_reset_out_reset),                                   //                   Nios2_reset_reset_bridge_in_reset.reset
		.JTAG_to_FPGA_Bridge_master_address                        (jtag_to_fpga_bridge_master_address),                                   //                          JTAG_to_FPGA_Bridge_master.address
		.JTAG_to_FPGA_Bridge_master_waitrequest                    (jtag_to_fpga_bridge_master_waitrequest),                               //                                                    .waitrequest
		.JTAG_to_FPGA_Bridge_master_byteenable                     (jtag_to_fpga_bridge_master_byteenable),                                //                                                    .byteenable
		.JTAG_to_FPGA_Bridge_master_read                           (jtag_to_fpga_bridge_master_read),                                      //                                                    .read
		.JTAG_to_FPGA_Bridge_master_readdata                       (jtag_to_fpga_bridge_master_readdata),                                  //                                                    .readdata
		.JTAG_to_FPGA_Bridge_master_readdatavalid                  (jtag_to_fpga_bridge_master_readdatavalid),                             //                                                    .readdatavalid
		.JTAG_to_FPGA_Bridge_master_write                          (jtag_to_fpga_bridge_master_write),                                     //                                                    .write
		.JTAG_to_FPGA_Bridge_master_writedata                      (jtag_to_fpga_bridge_master_writedata),                                 //                                                    .writedata
		.Nios2_data_master_address                                 (nios2_data_master_address),                                            //                                   Nios2_data_master.address
		.Nios2_data_master_waitrequest                             (nios2_data_master_waitrequest),                                        //                                                    .waitrequest
		.Nios2_data_master_byteenable                              (nios2_data_master_byteenable),                                         //                                                    .byteenable
		.Nios2_data_master_read                                    (nios2_data_master_read),                                               //                                                    .read
		.Nios2_data_master_readdata                                (nios2_data_master_readdata),                                           //                                                    .readdata
		.Nios2_data_master_write                                   (nios2_data_master_write),                                              //                                                    .write
		.Nios2_data_master_writedata                               (nios2_data_master_writedata),                                          //                                                    .writedata
		.Nios2_data_master_debugaccess                             (nios2_data_master_debugaccess),                                        //                                                    .debugaccess
		.Nios2_instruction_master_address                          (nios2_instruction_master_address),                                     //                            Nios2_instruction_master.address
		.Nios2_instruction_master_waitrequest                      (nios2_instruction_master_waitrequest),                                 //                                                    .waitrequest
		.Nios2_instruction_master_read                             (nios2_instruction_master_read),                                        //                                                    .read
		.Nios2_instruction_master_readdata                         (nios2_instruction_master_readdata),                                    //                                                    .readdata
		.VGA_Subsystem_pixel_dma_master_address                    (vga_subsystem_pixel_dma_master_address),                               //                      VGA_Subsystem_pixel_dma_master.address
		.VGA_Subsystem_pixel_dma_master_waitrequest                (vga_subsystem_pixel_dma_master_waitrequest),                           //                                                    .waitrequest
		.VGA_Subsystem_pixel_dma_master_read                       (vga_subsystem_pixel_dma_master_read),                                  //                                                    .read
		.VGA_Subsystem_pixel_dma_master_readdata                   (vga_subsystem_pixel_dma_master_readdata),                              //                                                    .readdata
		.VGA_Subsystem_pixel_dma_master_readdatavalid              (vga_subsystem_pixel_dma_master_readdatavalid),                         //                                                    .readdatavalid
		.VGA_Subsystem_pixel_dma_master_lock                       (vga_subsystem_pixel_dma_master_lock),                                  //                                                    .lock
		.Arduino_GPIO_s1_address                                   (mm_interconnect_0_arduino_gpio_s1_address),                            //                                     Arduino_GPIO_s1.address
		.Arduino_GPIO_s1_write                                     (mm_interconnect_0_arduino_gpio_s1_write),                              //                                                    .write
		.Arduino_GPIO_s1_readdata                                  (mm_interconnect_0_arduino_gpio_s1_readdata),                           //                                                    .readdata
		.Arduino_GPIO_s1_writedata                                 (mm_interconnect_0_arduino_gpio_s1_writedata),                          //                                                    .writedata
		.Arduino_GPIO_s1_chipselect                                (mm_interconnect_0_arduino_gpio_s1_chipselect),                         //                                                    .chipselect
		.Arduino_Reset_N_s1_address                                (mm_interconnect_0_arduino_reset_n_s1_address),                         //                                  Arduino_Reset_N_s1.address
		.Arduino_Reset_N_s1_write                                  (mm_interconnect_0_arduino_reset_n_s1_write),                           //                                                    .write
		.Arduino_Reset_N_s1_readdata                               (mm_interconnect_0_arduino_reset_n_s1_readdata),                        //                                                    .readdata
		.Arduino_Reset_N_s1_writedata                              (mm_interconnect_0_arduino_reset_n_s1_writedata),                       //                                                    .writedata
		.Arduino_Reset_N_s1_chipselect                             (mm_interconnect_0_arduino_reset_n_s1_chipselect),                      //                                                    .chipselect
		.HEX3_HEX0_s1_address                                      (mm_interconnect_0_hex3_hex0_s1_address),                               //                                        HEX3_HEX0_s1.address
		.HEX3_HEX0_s1_write                                        (mm_interconnect_0_hex3_hex0_s1_write),                                 //                                                    .write
		.HEX3_HEX0_s1_readdata                                     (mm_interconnect_0_hex3_hex0_s1_readdata),                              //                                                    .readdata
		.HEX3_HEX0_s1_writedata                                    (mm_interconnect_0_hex3_hex0_s1_writedata),                             //                                                    .writedata
		.HEX3_HEX0_s1_chipselect                                   (mm_interconnect_0_hex3_hex0_s1_chipselect),                            //                                                    .chipselect
		.HEX5_HEX4_s1_address                                      (mm_interconnect_0_hex5_hex4_s1_address),                               //                                        HEX5_HEX4_s1.address
		.HEX5_HEX4_s1_write                                        (mm_interconnect_0_hex5_hex4_s1_write),                                 //                                                    .write
		.HEX5_HEX4_s1_readdata                                     (mm_interconnect_0_hex5_hex4_s1_readdata),                              //                                                    .readdata
		.HEX5_HEX4_s1_writedata                                    (mm_interconnect_0_hex5_hex4_s1_writedata),                             //                                                    .writedata
		.HEX5_HEX4_s1_chipselect                                   (mm_interconnect_0_hex5_hex4_s1_chipselect),                            //                                                    .chipselect
		.Interval_Timer_s1_address                                 (mm_interconnect_0_interval_timer_s1_address),                          //                                   Interval_Timer_s1.address
		.Interval_Timer_s1_write                                   (mm_interconnect_0_interval_timer_s1_write),                            //                                                    .write
		.Interval_Timer_s1_readdata                                (mm_interconnect_0_interval_timer_s1_readdata),                         //                                                    .readdata
		.Interval_Timer_s1_writedata                               (mm_interconnect_0_interval_timer_s1_writedata),                        //                                                    .writedata
		.Interval_Timer_s1_chipselect                              (mm_interconnect_0_interval_timer_s1_chipselect),                       //                                                    .chipselect
		.Interval_Timer_2_s1_address                               (mm_interconnect_0_interval_timer_2_s1_address),                        //                                 Interval_Timer_2_s1.address
		.Interval_Timer_2_s1_write                                 (mm_interconnect_0_interval_timer_2_s1_write),                          //                                                    .write
		.Interval_Timer_2_s1_readdata                              (mm_interconnect_0_interval_timer_2_s1_readdata),                       //                                                    .readdata
		.Interval_Timer_2_s1_writedata                             (mm_interconnect_0_interval_timer_2_s1_writedata),                      //                                                    .writedata
		.Interval_Timer_2_s1_chipselect                            (mm_interconnect_0_interval_timer_2_s1_chipselect),                     //                                                    .chipselect
		.JTAG_UART_avalon_jtag_slave_address                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                //                         JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                  //                                                    .write
		.JTAG_UART_avalon_jtag_slave_read                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                   //                                                    .read
		.JTAG_UART_avalon_jtag_slave_readdata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),               //                                                    .readdata
		.JTAG_UART_avalon_jtag_slave_writedata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),              //                                                    .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),            //                                                    .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),             //                                                    .chipselect
		.LEDs_s1_address                                           (mm_interconnect_0_leds_s1_address),                                    //                                             LEDs_s1.address
		.LEDs_s1_write                                             (mm_interconnect_0_leds_s1_write),                                      //                                                    .write
		.LEDs_s1_readdata                                          (mm_interconnect_0_leds_s1_readdata),                                   //                                                    .readdata
		.LEDs_s1_writedata                                         (mm_interconnect_0_leds_s1_writedata),                                  //                                                    .writedata
		.LEDs_s1_chipselect                                        (mm_interconnect_0_leds_s1_chipselect),                                 //                                                    .chipselect
		.neopixel_0_avalon_slave_0_write                           (mm_interconnect_0_neopixel_0_avalon_slave_0_write),                    //                           neopixel_0_avalon_slave_0.write
		.neopixel_0_avalon_slave_0_writedata                       (mm_interconnect_0_neopixel_0_avalon_slave_0_writedata),                //                                                    .writedata
		.neopixel_0_avalon_slave_0_chipselect                      (mm_interconnect_0_neopixel_0_avalon_slave_0_chipselect),               //                                                    .chipselect
		.Nios2_debug_mem_slave_address                             (mm_interconnect_0_nios2_debug_mem_slave_address),                      //                               Nios2_debug_mem_slave.address
		.Nios2_debug_mem_slave_write                               (mm_interconnect_0_nios2_debug_mem_slave_write),                        //                                                    .write
		.Nios2_debug_mem_slave_read                                (mm_interconnect_0_nios2_debug_mem_slave_read),                         //                                                    .read
		.Nios2_debug_mem_slave_readdata                            (mm_interconnect_0_nios2_debug_mem_slave_readdata),                     //                                                    .readdata
		.Nios2_debug_mem_slave_writedata                           (mm_interconnect_0_nios2_debug_mem_slave_writedata),                    //                                                    .writedata
		.Nios2_debug_mem_slave_byteenable                          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),                   //                                                    .byteenable
		.Nios2_debug_mem_slave_waitrequest                         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),                  //                                                    .waitrequest
		.Nios2_debug_mem_slave_debugaccess                         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),                  //                                                    .debugaccess
		.Onchip_SRAM_s1_address                                    (mm_interconnect_0_onchip_sram_s1_address),                             //                                      Onchip_SRAM_s1.address
		.Onchip_SRAM_s1_write                                      (mm_interconnect_0_onchip_sram_s1_write),                               //                                                    .write
		.Onchip_SRAM_s1_readdata                                   (mm_interconnect_0_onchip_sram_s1_readdata),                            //                                                    .readdata
		.Onchip_SRAM_s1_writedata                                  (mm_interconnect_0_onchip_sram_s1_writedata),                           //                                                    .writedata
		.Onchip_SRAM_s1_byteenable                                 (mm_interconnect_0_onchip_sram_s1_byteenable),                          //                                                    .byteenable
		.Onchip_SRAM_s1_chipselect                                 (mm_interconnect_0_onchip_sram_s1_chipselect),                          //                                                    .chipselect
		.Onchip_SRAM_s1_clken                                      (mm_interconnect_0_onchip_sram_s1_clken),                               //                                                    .clken
		.Onchip_SRAM_s2_address                                    (mm_interconnect_0_onchip_sram_s2_address),                             //                                      Onchip_SRAM_s2.address
		.Onchip_SRAM_s2_write                                      (mm_interconnect_0_onchip_sram_s2_write),                               //                                                    .write
		.Onchip_SRAM_s2_readdata                                   (mm_interconnect_0_onchip_sram_s2_readdata),                            //                                                    .readdata
		.Onchip_SRAM_s2_writedata                                  (mm_interconnect_0_onchip_sram_s2_writedata),                           //                                                    .writedata
		.Onchip_SRAM_s2_byteenable                                 (mm_interconnect_0_onchip_sram_s2_byteenable),                          //                                                    .byteenable
		.Onchip_SRAM_s2_chipselect                                 (mm_interconnect_0_onchip_sram_s2_chipselect),                          //                                                    .chipselect
		.Onchip_SRAM_s2_clken                                      (mm_interconnect_0_onchip_sram_s2_clken),                               //                                                    .clken
		.Pushbuttons_s1_address                                    (mm_interconnect_0_pushbuttons_s1_address),                             //                                      Pushbuttons_s1.address
		.Pushbuttons_s1_write                                      (mm_interconnect_0_pushbuttons_s1_write),                               //                                                    .write
		.Pushbuttons_s1_readdata                                   (mm_interconnect_0_pushbuttons_s1_readdata),                            //                                                    .readdata
		.Pushbuttons_s1_writedata                                  (mm_interconnect_0_pushbuttons_s1_writedata),                           //                                                    .writedata
		.Pushbuttons_s1_chipselect                                 (mm_interconnect_0_pushbuttons_s1_chipselect),                          //                                                    .chipselect
		.SDRAM_s1_address                                          (mm_interconnect_0_sdram_s1_address),                                   //                                            SDRAM_s1.address
		.SDRAM_s1_write                                            (mm_interconnect_0_sdram_s1_write),                                     //                                                    .write
		.SDRAM_s1_read                                             (mm_interconnect_0_sdram_s1_read),                                      //                                                    .read
		.SDRAM_s1_readdata                                         (mm_interconnect_0_sdram_s1_readdata),                                  //                                                    .readdata
		.SDRAM_s1_writedata                                        (mm_interconnect_0_sdram_s1_writedata),                                 //                                                    .writedata
		.SDRAM_s1_byteenable                                       (mm_interconnect_0_sdram_s1_byteenable),                                //                                                    .byteenable
		.SDRAM_s1_readdatavalid                                    (mm_interconnect_0_sdram_s1_readdatavalid),                             //                                                    .readdatavalid
		.SDRAM_s1_waitrequest                                      (mm_interconnect_0_sdram_s1_waitrequest),                               //                                                    .waitrequest
		.SDRAM_s1_chipselect                                       (mm_interconnect_0_sdram_s1_chipselect),                                //                                                    .chipselect
		.servo_0_avalon_slave_0_write                              (mm_interconnect_0_servo_0_avalon_slave_0_write),                       //                              servo_0_avalon_slave_0.write
		.servo_0_avalon_slave_0_writedata                          (mm_interconnect_0_servo_0_avalon_slave_0_writedata),                   //                                                    .writedata
		.servo_0_avalon_slave_0_chipselect                         (mm_interconnect_0_servo_0_avalon_slave_0_chipselect),                  //                                                    .chipselect
		.Slider_Switches_s1_address                                (mm_interconnect_0_slider_switches_s1_address),                         //                                  Slider_Switches_s1.address
		.Slider_Switches_s1_readdata                               (mm_interconnect_0_slider_switches_s1_readdata),                        //                                                    .readdata
		.SysID_control_slave_address                               (mm_interconnect_0_sysid_control_slave_address),                        //                                 SysID_control_slave.address
		.SysID_control_slave_readdata                              (mm_interconnect_0_sysid_control_slave_readdata),                       //                                                    .readdata
		.telemetre_0_avalon_slave_0_read                           (mm_interconnect_0_telemetre_0_avalon_slave_0_read),                    //                          telemetre_0_avalon_slave_0.read
		.telemetre_0_avalon_slave_0_readdata                       (mm_interconnect_0_telemetre_0_avalon_slave_0_readdata),                //                                                    .readdata
		.telemetre_0_avalon_slave_0_chipselect                     (mm_interconnect_0_telemetre_0_avalon_slave_0_chipselect),              //                                                    .chipselect
		.uart_0_avalon_slave_0_write                               (mm_interconnect_0_uart_0_avalon_slave_0_write),                        //                               uart_0_avalon_slave_0.write
		.uart_0_avalon_slave_0_read                                (mm_interconnect_0_uart_0_avalon_slave_0_read),                         //                                                    .read
		.uart_0_avalon_slave_0_readdata                            (mm_interconnect_0_uart_0_avalon_slave_0_readdata),                     //                                                    .readdata
		.uart_0_avalon_slave_0_writedata                           (mm_interconnect_0_uart_0_avalon_slave_0_writedata),                    //                                                    .writedata
		.VGA_Subsystem_char_buffer_control_slave_address           (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address),    //             VGA_Subsystem_char_buffer_control_slave.address
		.VGA_Subsystem_char_buffer_control_slave_write             (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write),      //                                                    .write
		.VGA_Subsystem_char_buffer_control_slave_read              (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read),       //                                                    .read
		.VGA_Subsystem_char_buffer_control_slave_readdata          (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata),   //                                                    .readdata
		.VGA_Subsystem_char_buffer_control_slave_writedata         (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata),  //                                                    .writedata
		.VGA_Subsystem_char_buffer_control_slave_byteenable        (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable), //                                                    .byteenable
		.VGA_Subsystem_char_buffer_slave_address                   (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),            //                     VGA_Subsystem_char_buffer_slave.address
		.VGA_Subsystem_char_buffer_slave_write                     (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),              //                                                    .write
		.VGA_Subsystem_char_buffer_slave_readdata                  (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),           //                                                    .readdata
		.VGA_Subsystem_char_buffer_slave_writedata                 (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),          //                                                    .writedata
		.VGA_Subsystem_char_buffer_slave_byteenable                (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),         //                                                    .byteenable
		.VGA_Subsystem_char_buffer_slave_chipselect                (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect),         //                                                    .chipselect
		.VGA_Subsystem_char_buffer_slave_clken                     (mm_interconnect_0_vga_subsystem_char_buffer_slave_clken),              //                                                    .clken
		.VGA_Subsystem_pixel_dma_control_slave_address             (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),      //               VGA_Subsystem_pixel_dma_control_slave.address
		.VGA_Subsystem_pixel_dma_control_slave_write               (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),        //                                                    .write
		.VGA_Subsystem_pixel_dma_control_slave_read                (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),         //                                                    .read
		.VGA_Subsystem_pixel_dma_control_slave_readdata            (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),     //                                                    .readdata
		.VGA_Subsystem_pixel_dma_control_slave_writedata           (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),    //                                                    .writedata
		.VGA_Subsystem_pixel_dma_control_slave_byteenable          (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable),   //                                                    .byteenable
		.VGA_Subsystem_rgb_slave_read                              (mm_interconnect_0_vga_subsystem_rgb_slave_read),                       //                             VGA_Subsystem_rgb_slave.read
		.VGA_Subsystem_rgb_slave_readdata                          (mm_interconnect_0_vga_subsystem_rgb_slave_readdata)                    //                                                    .readdata
	);

	Computer_System_irq_mapper irq_mapper (
		.clk           (system_pll_sys_clk_clk),             //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (system_pll_reset_source_reset),      // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_debug_reset_request_reset),    // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
